----------------------------------------------------------
--Description: top entity with instance of the pipe levels
--and registers among them
--the processor has to exchange data with the external
--data and instruction memories
----------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity RISC_V is
    port(
        RISC_V_IN_RST_N         : in std_logic;
        RISC_V_IN_CLK           : in std_logic;
        RISC_V_IN_INSTR         : in std_logic_vector(31 downto 0);        --instruction read from the code memory
        RISC_V_IN_RD_DATA       : in std_logic_vector(31 downto 0);        --data read from data memory
        RISC_V_OUT_PC           : out std_logic_vector(31 downto 0);       --program counter
        RISC_V_OUT_WR_DATA      : out std_logic_vector(31 downto 0);       --data written in the data memory
        RISC_V_OUT_WR_ADD       : out std_logic_vector(31 downto 0);       --address for the write in the data memory
        RISC_V_OUT_MEMWRITE     : out std_logic;                           --control signal of the data memory
        RISC_V_OUT_MEMREAD      : out std_logic                            --control signal of the data memory
    );
end entity;

architecture structural of RISC_V is
    component instr_fetch is
        port (
            INSTR_FETCH_IN_PC_WRBRANCH: in std_logic_vector(31 downto 0);     --address to take in case of wrong branch
            INSTR_FETCH_IN_BRANCH    : in std_logic;                          --signal to detect if a jump has to be performed
            INSTR_FETCH_IN_RST_N     : in std_logic;                          --reset for PC
            INSTR_FETCH_IN_CLK       : in std_logic;                          --clock for PC
            INSTR_FETCH_IN_PC_EN     : in std_logic;                          --pc register enable
            INSTR_FETCH_IN_WRONGPRED : in std_logic;                          --signal to understand if the branch prediction was wrong
            INSTR_FETCH_IN_WADD_PBTAB: in std_logic_vector(31 downto 0);       --write address of the PB table
            INSTR_FETCH_IN_INSTR     : in std_logic_vector(31 downto 0);      --instruction from memory
            INSTR_FETCH_OUT_INSTR    : out std_logic_vector(31 downto 0);     --instruction for decode stage
            INSTR_FETCH_OUT_ADDR     : out std_logic_vector(31 downto 0);     --address for memory
            INSTR_FETCH_OUT_BRANCHPRED: out std_logic                         --branch prediction bit read from the BPtable
        );
    end component;
    signal pc_branch_from_mem_stage, instruction_from_fetch_stage, pc_from_fetch_stage   : std_logic_vector(31 downto 0);
    signal pcsrc_from_mem_stage,branch_pred_from_fetch_stage                             : std_logic;

    component DECODE_STAGE is
        port(

            DEC_STAGE_IN_INSTR : in std_logic_vector(31 downto 0); --instruction fecthed from IM
            DEC_STAGE_IN_PC    : in std_logic_vector(31 downto 0); --program counter
            DEC_STAGE_OUT_JAL        : out std_logic;                     --signal to jump for jar operation
            DEC_STAGE_OUT_BRANCH     : out std_logic;                     --signal to dected if a branch is fetched
            DEC_STAGE_OUT_MEMREAD    : out std_logic;                     --control signal for the data memory
            DEC_STAGE_OUT_MEMWRITE   : out std_logic;                     --control signal for the data memory
            DEC_STAGE_OUT_MEMTOREG   : out std_logic;                     --control signal for the data memory
            DEC_STAGE_OUT_REGWRITE   : out std_logic;                     --signal to write in the register file generated by CU
            DEC_STAGE_OUT_ALUSRC1    : out std_logic;                     --selection signal mux at the input of the ALU
            DEC_STAGE_OUT_ALUSRC2    : out std_logic_vector(1 downto 0);  --selection signal mux at the input of the ALU
            DEC_STAGE_OUT_ALURES     : out std_logic;                     --selection signal mux at the output of the ALU
            DEC_STAGE_OUT_ALUOP      : out std_logic_vector(1 downto 0);  --output CU for the ALUControl

            DEC_STAGE_IN_CLK       : in std_logic;                      -- clock of the register file

            DEC_STAGE_IN_REGWRITE  : in std_logic;                      --signal to write in the register file from WB stage
            DEC_STAGE_IN_WRITEADD  : in std_logic_vector(4 downto 0);   --write address
            DEC_STAGE_IN_WRITEDATA : in std_logic_vector(31 downto 0);  --write data

            DEC_STAGE_OUT_READDATA1 : out std_logic_vector(31 downto 0); --first output register file
            DEC_STAGE_OUT_READDATA2 : out std_logic_vector(31 downto 0); --second output register file

            DEC_STAGE_OUT_IMM : out std_logic_vector(31 downto 0);  --output immediate generation unit

            --hazard detection useful signals
            DEC_STAGE_IN_MEMREAD_ID_EX : in std_logic;
            DEC_STAGE_IN_RD_ID_EX      : in std_logic_vector(4 downto 0);
            DEC_OUT_PC_EN              : out std_logic;
            DEC_OUT_IF_ID_LOAD         : out std_logic;

            DEC_STAGE_OUT_FUNC4 : out std_logic_vector(3 downto 0); --field used by alu control
            DEC_STAGE_OUT_RS1   : out std_logic_vector(4 downto 0); --source1 register field
            DEC_STAGE_OUT_RS2   : out std_logic_vector(4 downto 0); --source2 register field
            DEC_STAGE_OUT_RD    : out std_logic_vector(4 downto 0); --destination register field
            DEC_STAGE_OUT_PC    : out std_logic_vector(31 downto 0) --program counter

        );
      end component;

    signal branch_from_decode_stage, jal_from_decode_stage, memread_from_decode_stage, memwrite_from_decode_stage, memtoreg_from_decode_stage  : std_logic;
    signal regwrite_from_decode_stage, alusrc1_from_decode_stage, alures_from_decode_stage                                                     : std_logic;
    signal alusrc2_from_decode_stage, aluop_from_decode_stage                                                                                  : std_logic_vector (1 downto 0);
    signal read_data1_from_decode_stage, read_data2_from_decode_stage, immediate_from_decode_stage, pc_from_decode_stage                       : std_logic_vector (31 downto 0);
    signal func4_from_decode_stage                                                                                                             : std_logic_vector(3 downto 0);
    signal rd_from_decode_stage, rs1_from_decode_stage, rs2_from_decode_stage                                                                  : std_logic_vector(4 downto 0);
    signal pc_en_from_dec_to_fetch                                                                                                             : std_logic;    --program counter enable
    signal if_dec_reg_en                                                                                                                       : std_logic;    --enable of IF/DEC pipe register

    component EXECUTION_STAGE is
        port (
            EXEC_STAGE_IN_IMM_GEN         : in std_logic_vector(31 downto 0); --output immediate generation unit
            EXEC_STAGE_IN_PC              : in std_logic_vector(31 downto 0); --program counter
            EXEC_STAGE_IN_DATA1           : in std_logic_vector(31 downto 0); --first output register file
            EXEC_STAGE_IN_DATA2           : in std_logic_vector(31 downto 0); --second output register file
            EXEC_STAGE_IN_SHORT_BYPASS    : in std_logic_vector(31 downto 0); --prior ALU result (1 delay)
            EXEC_STAGE_IN_LONG_BYPASS     : in std_logic_vector(31 downto 0); --earlier ALU result (2 delay) or data memory value (1 delay)
            EXEC_STAGE_IN_ALUOP           : in std_logic_vector(1 downto 0);  --output CU for the ALUControl
            EXEC_STAGE_IN_FUNC4           : in std_logic_vector(3 downto 0);  --field used BY alu control
            EXEC_STAGE_IN_ALUSRC1         : in std_logic;                     -- selection signal mux at the input of the ALU
            EXEC_STAGE_IN_ALUSRC2         : in std_logic_vector(1 downto 0);  -- selection signal mux at the input of the ALU
            EXEC_STAGE_IN_ALURES          : in std_logic;                     -- selection signal mux at the output of the ALU
            EXEC_STAGE_IN_MEMREAD         : in std_logic;                     --control signal for the data memory
            EXEC_STAGE_IN_MEMWRITE        : in std_logic;                     --control signal for the data memory
            EXEC_STAGE_IN_MEMTOREG        : in std_logic;                     --control signal for the data memory
            EXEC_STAGE_IN_BRANCH          : in std_logic;                     --signal to dected if a BEQ is fetched
            EXEC_STAGE_IN_JAL             : in std_logic;                     --signal to jump for JAL op
            EXEC_STAGE_IN_REGWRITE        : in std_logic;                     --signal to write in the register file
            EXEC_STAGE_IN_REGWRITE_EX_MEM : in std_logic;                     --signal to write in the register file from ex_mem stage
            EXEC_STAGE_IN_REGWRITE_MEM_WB : in std_logic;                     --signal to write in the register file from mem_wb stage
            EXEC_STAGE_IN_SR1             : in std_logic_vector(4 downto 0);  --address of the source1 register
            EXEC_STAGE_IN_SR2             : in std_logic_vector(4 downto 0);  --address of the source2 register
            EXEC_STAGE_IN_RD              : in std_logic_vector(4 downto 0);  --address of the destination register
            EXEC_STAGE_IN_RD_EX_MEM       : in std_logic_vector(4 downto 0);  --address of the destination register from ex_mem stage
            EXEC_STAGE_IN_RD_MEM_WB       : in std_logic_vector(4 downto 0);  --address of the destination register from mem_wb stage
            EXEC_STAGE_OUT_ALU            : out std_logic_vector(31 downto 0);-- ALU output
            EXEC_STAGE_OUT_PC_BRANCH      : out std_logic_vector(31 downto 0);--PC evaluated in case of branch
            EXEC_STAGE_OUT_ZERO_FLAG      : out std_logic;                    --zero flag of the ALU
            EXEC_STAGE_OUT_SRC2           : out std_logic_vector(31 downto 0);--second output register file
            EXEC_STAGE_OUT_RD             : out std_logic_vector(4 downto 0); --address of the destination register
            EXEC_STAGE_OUT_MEMREAD        : out std_logic;                    --control signal for the data memory
            EXEC_STAGE_OUT_MEMWRITE       : out std_logic;                    --control signal for the data memory
            EXEC_STAGE_OUT_MEMTOREG       : out std_logic;                    --control signal for the data memory
            EXEC_STAGE_OUT_BRANCH         : out std_logic;                    --signal to dected if a BEQ is fetched
            EXEC_STAGE_OUT_JAL            : out std_logic;                    --signal to jump for JAL op
            EXEC_STAGE_OUT_REGWRITE       : out std_logic;                     --signal to write in the register file
            EXEC_STAGE_IN_CLK             : in std_logic;                     --used by CHDU flip-flops
            EXEC_STAGE_IN_FLUSH           : in std_logic;                     --signal to flush the pipe
            EXEC_STAGE_IN_BRANCHPRED      : in std_logic;                     --signal to know if a jump is predicted or not
            EXEC_STAGE_OUT_BRANCHPRED     : out std_logic                     --signal to know if a jump is predicted or not
        );
    end component;

    signal zero_flag_from_execution_stage, branch_from_execution_stage, jal_from_execution_stage, memwrite_from_execution_stage    : std_logic;
    signal memread_from_execution_stage, regwrite_from_execution_stage, memtoreg_from_execution_stage                              : std_logic;
    signal branchpred_from_execution_stage                                                                                         : std_logic;
    signal pc_branch_from_execution_stage, write_data_from_execution_stage, alu_res_from_execution_stage                           : std_logic_vector (31 downto 0);
    signal rd_from_execution_stage                                                                                                 : std_logic_vector (4 downto 0);


    component memory_stage is
        port (
            MEM_STAGE_IN_ZERO_F      : in std_logic;                        --zero flag from execution stage
            MEM_STAGE_IN_BRANCH      : in std_logic;                        --control branch from EU
            MEM_STAGE_IN_JAL         : in std_logic;                        --jump for jal from EU
            MEM_STAGE_IN_MEMWRITE    : in std_logic;                        --control write mem from EU
            MEM_STAGE_IN_MEMREAD     : in std_logic;                        --control read mem from EU
            MEM_STAGE_IN_REGWRITE    : in std_logic;                        --control write RF from EU
            MEM_STAGE_IN_MEMTOREG    : in std_logic;                        --control to decide what to write back in the register file
            MEM_STAGE_IN_ALU_RES     : in std_logic_vector(31 downto 0);    --result of the alu from the exec stage
            MEM_STAGE_IN_WR_DATA     : in std_logic_vector(31 downto 0);    --data to write in memory from execution stage
            MEM_STAGE_IN_RD_DATA     : in std_logic_vector(31 downto 0);    --data read from data memory
            MEM_STAGE_IN_PC_BRANCH   : in std_logic_vector(31 downto 0);    --address to jump for fetch stage
            MEM_STAGE_IN_RD          : in std_logic_vector(4 downto 0);     --destination register for the write back
            MEM_STAGE_IN_BRANCHPRED  : in std_logic;                        --signal with the branch prediction of the PBtable
            MEM_STAGE_OUT_BRANCH     : out std_logic;                       --control to decide if jump or not, for fetch stage
            MEM_STAGE_OUT_MEMWRITE   : out std_logic;                       --control write for data memory
            MEM_STAGE_OUT_MEMREAD    : out std_logic;                       --control read for data memory
            MEM_STAGE_OUT_REGWRITE   : out std_logic;                       --control write for RF
            MEM_STAGE_OUT_MEMTOREG   : out std_logic;                       --control to decide what to write back in the register file
            MEM_STAGE_OUT_ALU_RES    : out std_logic_vector(31 downto 0);   --result of the alu from the exec stage
            MEM_STAGE_OUT_WR_DATA    : out std_logic_vector(31 downto 0);   --data that has to written in the data memory
            MEM_STAGE_OUT_RD_DATA    : out std_logic_vector(31 downto 0);    --data read from the data memory
            MEM_STAGE_OUT_PC_WRBRANCH: out std_logic_vector(31 downto 0);   --address to jump in case of wrong branch prediction
            MEM_STAGE_OUT_RD         : out std_logic_vector(4 downto 0);    --destination register for the write back
            MEM_STAGE_OUT_WRONGPRED  : out std_logic                        --signal to understand if the branch prediction was wrong
        );
    end component;

    signal zero_flag_to_mem_stage, branch_to_mem_stage, jal_to_mem_stage, regwrite_from_mem_stage,  memwrite_to_mem_stage       : std_logic;
    signal memread_to_mem_stage, regwrite_to_mem_stage, memtoreg_to_mem_stage, memtoreg_from_mem_stage, wrongpred_from_mem_stage: std_logic;
    signal alu_res_to_mem_stage, alu_res_from_mem_stage, write_data_to_mem_stage, pc_wrbranch_to_mem_stage                      : std_logic_vector (31 downto 0);
    signal pc_wrbranch_from_mem_stage, rd_data_from_mem_stage, pc_from_mem_stage, pc_branch_to_mem_stage                        : std_logic_vector (31 downto 0);
    signal rd_to_mem_stage, rd_from_mem_stage                                                                                   : std_logic_vector (4 downto 0);

    component REGISTER_NBIT is
        generic (N_g:integer:=8);
        port (
            REGISTER_IN_RST_N  : in std_logic;
            REGISTER_IN_CLK    : in std_logic;
            REGISTER_IN_EN     : in std_logic;
            REGISTER_IN_D      : in std_logic_vector(N_g-1 downto 0);
            REGISTER_OUT_Q     : out std_logic_vector(N_g-1 downto 0)
        );
    end component;
    signal reg_IF_ID_in, reg_IF_ID_out   : std_logic_vector (64 downto 0);
    signal reg_EX_MEM_in, reg_EX_MEM_out : std_logic_vector (140 downto 0);
    signal reg_MEM_WB_in, reg_MEM_WB_out : std_logic_vector (70 downto 0);
    signal reg_ID_EX_in, reg_ID_EX_out   : std_logic_vector (159 downto 0);

    component MUX2TO1 is
        generic(N_g: integer:=4);
        port(
            MUX_IN_D0   : IN std_logic_vector (N_g-1 downto 0);
            MUX_IN_D1   : IN std_logic_vector (N_g-1 downto 0);
            MUX_IN_SEL  : IN std_logic;
            MUX_OUT     : OUT std_logic_vector (N_g-1 downto 0)
        );
    end component;

    signal rd_from_wb_stage         : std_logic_vector(4 downto 0);
    signal regwrite_from_wb_stage   : std_logic;
    signal output_from_wb_stage     : std_logic_vector(31 downto 0);


    begin

        i_fetch_stage: instr_fetch
            port map(
            INSTR_FETCH_IN_PC_WRBRANCH=> pc_wrbranch_from_mem_stage,
            INSTR_FETCH_IN_BRANCH    => pcsrc_from_mem_stage,
            INSTR_FETCH_IN_RST_N     => RISC_V_IN_RST_N,
            INSTR_FETCH_IN_CLK       => RISC_V_IN_CLK,
            INSTR_FETCH_IN_PC_EN     => pc_en_from_dec_to_fetch,
            INSTR_FETCH_IN_WRONGPRED => wrongpred_from_mem_stage,
            INSTR_FETCH_IN_WADD_PBTAB=> pc_from_mem_stage,
            INSTR_FETCH_IN_INSTR     => RISC_V_IN_INSTR,
            INSTR_FETCH_OUT_INSTR    => instruction_from_fetch_stage,
            INSTR_FETCH_OUT_ADDR     => pc_from_fetch_stage,
            INSTR_FETCH_OUT_BRANCHPRED=> branch_pred_from_fetch_stage
            );
        RISC_V_OUT_PC  <=  pc_from_fetch_stage;

        reg_IF_ID_in   <= branch_pred_from_fetch_stage & instruction_from_fetch_stage & pc_from_fetch_stage;
        --dimension: PC+ instruction
        i_reg_IF_ID: REGISTER_NBIT
            generic map (N_g=> 65)
            port map (
                REGISTER_IN_RST_N  => RISC_V_IN_RST_N,
                REGISTER_IN_CLK    => RISC_V_IN_CLK,
                REGISTER_IN_EN     => if_dec_reg_en,
                REGISTER_IN_D      => reg_IF_ID_in,
                REGISTER_OUT_Q     => reg_IF_ID_out
            );

        i_decode_stage: DECODE_STAGE
            port map(
                DEC_STAGE_IN_INSTR      => reg_IF_ID_out(63 downto 32),
                DEC_STAGE_IN_PC         => reg_IF_ID_out(31 downto 0),
                DEC_STAGE_OUT_JAL       => jal_from_decode_stage,
                DEC_STAGE_OUT_BRANCH    => branch_from_decode_stage,
                DEC_STAGE_OUT_MEMREAD   => memread_from_decode_stage,
                DEC_STAGE_OUT_MEMWRITE  => memwrite_from_decode_stage,
                DEC_STAGE_OUT_MEMTOREG  => memtoreg_from_decode_stage,
                DEC_STAGE_OUT_REGWRITE  => regwrite_from_decode_stage,
                DEC_STAGE_OUT_ALUSRC1   => alusrc1_from_decode_stage,
                DEC_STAGE_OUT_ALUSRC2   => alusrc2_from_decode_stage,
                DEC_STAGE_OUT_ALURES    => alures_from_decode_stage,
                DEC_STAGE_OUT_ALUOP     => aluop_from_decode_stage,
                DEC_STAGE_IN_CLK        => RISC_V_IN_CLK,
                DEC_STAGE_IN_REGWRITE      => regwrite_from_wb_stage,
                DEC_STAGE_IN_WRITEADD      => rd_from_wb_stage,
                DEC_STAGE_IN_WRITEDATA     => output_from_wb_stage,
                DEC_STAGE_OUT_READDATA1    => read_data1_from_decode_stage,
                DEC_STAGE_OUT_READDATA2    => read_data2_from_decode_stage,
                DEC_STAGE_OUT_IMM          => immediate_from_decode_stage,
                DEC_STAGE_IN_MEMREAD_ID_EX => memread_from_execution_stage,
                DEC_STAGE_IN_RD_ID_EX      => rd_from_execution_stage,
                DEC_OUT_PC_EN              => pc_en_from_dec_to_fetch,
                DEC_OUT_IF_ID_LOAD         => if_dec_reg_en,
                DEC_STAGE_OUT_FUNC4     => func4_from_decode_stage,
                DEC_STAGE_OUT_RS1       => rs1_from_decode_stage,
                DEC_STAGE_OUT_RS2       => rs2_from_decode_stage,
                DEC_STAGE_OUT_RD        => rd_from_decode_stage,
                DEC_STAGE_OUT_PC        => pc_from_decode_stage

            );

        reg_ID_EX_in   <= ( reg_IF_ID_out(64) & rs1_from_decode_stage & rs2_from_decode_stage & jal_from_decode_stage & branch_from_decode_stage & memread_from_decode_stage & memwrite_from_decode_stage & memtoreg_from_decode_stage
                            & regwrite_from_decode_stage & alusrc1_from_decode_stage & alusrc2_from_decode_stage & alures_from_decode_stage
                            & aluop_from_decode_stage & read_data1_from_decode_stage & read_data2_from_decode_stage & immediate_from_decode_stage &
                            func4_from_decode_stage & rd_from_decode_stage & pc_from_decode_stage);

        i_reg_ID_EX: REGISTER_NBIT
            generic map (N_g=> 160)
            port map (
                REGISTER_IN_RST_N  => RISC_V_IN_RST_N,
                REGISTER_IN_CLK    => RISC_V_IN_CLK,
                REGISTER_IN_EN     => '1',
                REGISTER_IN_D      => reg_ID_EX_in,
                REGISTER_OUT_Q     => reg_ID_EX_out
            );

        i_execution_stage: EXECUTION_STAGE
            port map(
                EXEC_STAGE_IN_IMM_GEN         => reg_ID_EX_out(72 downto 41),
                EXEC_STAGE_IN_PC              => reg_ID_EX_out(31 downto 0),
                EXEC_STAGE_IN_DATA1           => reg_ID_EX_out(136 downto 105),
                EXEC_STAGE_IN_DATA2           => reg_ID_EX_out(104 downto 73),
                EXEC_STAGE_IN_SHORT_BYPASS    => alu_res_to_mem_stage,
                EXEC_STAGE_IN_LONG_BYPASS     => output_from_wb_stage,
                EXEC_STAGE_IN_ALUOP           => reg_ID_EX_out(138 downto 137),
                EXEC_STAGE_IN_FUNC4           => reg_ID_EX_out(40 downto 37),
                EXEC_STAGE_IN_ALUSRC1         => reg_ID_EX_out(142),
                EXEC_STAGE_IN_ALUSRC2         => reg_ID_EX_out(141 downto 140),
                EXEC_STAGE_IN_ALURES          => reg_ID_EX_out(139),
                EXEC_STAGE_IN_MEMREAD         => reg_ID_EX_out(146),
                EXEC_STAGE_IN_MEMWRITE        => reg_ID_EX_out(145),
                EXEC_STAGE_IN_MEMTOREG        => reg_ID_EX_out(144),
                EXEC_STAGE_IN_BRANCH          => reg_ID_EX_out(147),
                EXEC_STAGE_IN_JAL             => reg_ID_EX_out(148),
                EXEC_STAGE_IN_REGWRITE        => reg_ID_EX_out(143),
                EXEC_STAGE_IN_REGWRITE_EX_MEM => regwrite_from_mem_stage,
                EXEC_STAGE_IN_REGWRITE_MEM_WB => regwrite_from_wb_stage,
                EXEC_STAGE_IN_SR1             => reg_ID_EX_out(158 downto 154),
                EXEC_STAGE_IN_SR2             => reg_ID_EX_out(153 downto 149),
                EXEC_STAGE_IN_RD              => reg_ID_EX_out(36 downto 32),
                EXEC_STAGE_IN_RD_EX_MEM       => rd_to_mem_stage,
                EXEC_STAGE_IN_RD_MEM_WB       => rd_from_wb_stage,
                EXEC_STAGE_OUT_ALU            => alu_res_from_execution_stage,
                EXEC_STAGE_OUT_PC_BRANCH      => pc_branch_from_execution_stage,
                EXEC_STAGE_OUT_ZERO_FLAG      => zero_flag_from_execution_stage,
                EXEC_STAGE_OUT_SRC2           => write_data_from_execution_stage,
                EXEC_STAGE_OUT_RD             => rd_from_execution_stage,
                EXEC_STAGE_OUT_MEMREAD        => memread_from_execution_stage,
                EXEC_STAGE_OUT_MEMWRITE       => memwrite_from_execution_stage,
                EXEC_STAGE_OUT_MEMTOREG       => memtoreg_from_execution_stage,
                EXEC_STAGE_OUT_BRANCH         => branch_from_execution_stage,
                EXEC_STAGE_OUT_JAL            => jal_from_execution_stage,
                EXEC_STAGE_OUT_REGWRITE       => regwrite_from_execution_stage,
                EXEC_STAGE_IN_CLK             => RISC_V_IN_CLK,
                EXEC_STAGE_IN_FLUSH           => wrongpred_from_mem_stage,
                EXEC_STAGE_IN_BRANCHPRED      => reg_ID_EX_out(159),
                EXEC_STAGE_OUT_BRANCHPRED     => branchpred_from_execution_stage
            );

            reg_EX_MEM_in <= (reg_ID_EX_out(31 downto 0) & branchpred_from_execution_stage & jal_from_execution_stage & zero_flag_from_execution_stage & branch_from_execution_stage & memwrite_from_execution_stage & memread_from_execution_stage
                            & regwrite_from_execution_stage & memtoreg_from_execution_stage & alu_res_from_execution_stage &
                            write_data_from_execution_stage & pc_branch_from_execution_stage & rd_from_execution_stage);
            --dimension: 3 control signals for the memory+zero flag+branch control+memtoreg control+ alu_re (32 bit) + write_data(32 bit)+pc_branch(32 bit)+ rd(5 bit)
            i_reg_EX_MEM: REGISTER_NBIT
                generic map (N_g=> 141)
                port map (
                    REGISTER_IN_RST_N  => RISC_V_IN_RST_N,
                    REGISTER_IN_CLK    => RISC_V_IN_CLK,
                    REGISTER_IN_EN     => '1',
                    REGISTER_IN_D      => reg_EX_MEM_in,
                    REGISTER_OUT_Q     => reg_EX_MEM_out
                );
            rd_to_mem_stage         <= reg_EX_MEM_out(4 downto 0);
            pc_branch_to_mem_stage  <= reg_EX_MEM_out(36 downto 5);
            write_data_to_mem_stage <= reg_EX_MEM_out(68 downto 37);
            alu_res_to_mem_stage    <= reg_EX_MEM_out(100 downto 69);
            memtoreg_to_mem_stage   <= reg_EX_MEM_out(101);
            regwrite_to_mem_stage   <= reg_EX_MEM_out(102);
            memread_to_mem_stage    <= reg_EX_MEM_out(103);
            memwrite_to_mem_stage   <= reg_EX_MEM_out(104);
            branch_to_mem_stage     <= reg_EX_MEM_out(105);
            zero_flag_to_mem_stage  <= reg_EX_MEM_out(106);
            jal_to_mem_stage        <= reg_EX_MEM_out(107);
            pc_from_mem_stage       <= reg_EX_MEM_out(140 downto 109);

            i_memory_stage: memory_stage
                port map(
                MEM_STAGE_IN_ZERO_F      => zero_flag_to_mem_stage,
                MEM_STAGE_IN_BRANCH      => branch_to_mem_stage,
                MEM_STAGE_IN_JAL         => jal_to_mem_stage,
                MEM_STAGE_IN_MEMWRITE    => memwrite_to_mem_stage,
                MEM_STAGE_IN_MEMREAD     => memread_to_mem_stage,
                MEM_STAGE_IN_REGWRITE    => regwrite_to_mem_stage,
                MEM_STAGE_IN_MEMTOREG    => memtoreg_to_mem_stage,
                MEM_STAGE_IN_ALU_RES     => alu_res_to_mem_stage,
                MEM_STAGE_IN_WR_DATA     => write_data_to_mem_stage,
                MEM_STAGE_IN_RD_DATA     => RISC_V_IN_RD_DATA,
                MEM_STAGE_IN_PC_BRANCH   => pc_branch_to_mem_stage,
                MEM_STAGE_IN_RD          => rd_to_mem_stage,
                MEM_STAGE_IN_BRANCHPRED  => reg_EX_MEM_out(108),
                MEM_STAGE_OUT_BRANCH     => pcsrc_from_mem_stage,
                MEM_STAGE_OUT_MEMWRITE   => RISC_V_OUT_MEMWRITE,
                MEM_STAGE_OUT_MEMREAD    => RISC_V_OUT_MEMREAD,
                MEM_STAGE_OUT_REGWRITE   => regwrite_from_mem_stage,
                MEM_STAGE_OUT_MEMTOREG   => memtoreg_from_mem_stage,
                MEM_STAGE_OUT_ALU_RES    => alu_res_from_mem_stage,
                MEM_STAGE_OUT_WR_DATA    => RISC_V_OUT_WR_DATA,
                MEM_STAGE_OUT_RD_DATA    => rd_data_from_mem_stage,
                MEM_STAGE_OUT_PC_WRBRANCH=> pc_wrbranch_from_mem_stage,
                MEM_STAGE_OUT_RD         => rd_from_mem_stage,
                MEM_STAGE_OUT_WRONGPRED  => wrongpred_from_mem_stage
                );

            RISC_V_OUT_WR_ADD <= alu_res_from_mem_stage;

            reg_MEM_WB_in <= (regwrite_from_mem_stage & memtoreg_from_mem_stage & alu_res_from_mem_stage
                                & rd_data_from_mem_stage & rd_from_mem_stage );
            i_reg_MEM_WB: REGISTER_NBIT
                generic map (N_g=> 71)
                port map (
                    REGISTER_IN_RST_N  => RISC_V_IN_RST_N,
                    REGISTER_IN_CLK    => RISC_V_IN_CLK,
                    REGISTER_IN_EN     => '1',
                    REGISTER_IN_D      => reg_MEM_WB_in,
                    REGISTER_OUT_Q     => reg_MEM_WB_out
                );

            rd_from_wb_stage         <= reg_MEM_WB_out(4 downto 0);
            regwrite_from_wb_stage   <= reg_MEM_WB_out(70);

            i_final_mux: MUX2TO1
                generic map(N_g=> 32)
                port map(
                    MUX_IN_D0   => reg_MEM_WB_out(68 downto 37),
                    MUX_IN_D1   => reg_MEM_WB_out(36 downto 5),
                    MUX_IN_SEL  => reg_MEM_WB_out(69),
                    MUX_OUT     => output_from_wb_stage
                );
end architecture;
