C:/software/dk/nangate45/lef/NangateOpenCellLibrary.lef